class scoreboard;
	mailbox scb_mbx;
