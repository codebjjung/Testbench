class Packet;
	rand bit [3:0] a;
	rand bit [3:0] b;
	bit [7:0] y;
endclass
