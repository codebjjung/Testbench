class Packet;
   rand bit [31:0] paddr;
   rand bit [31:0] pwdata;
   bit pwrite;
   bit psel;
   bit penable;
   bit [3:0] pstrb;
   bit prdata;
endclass
