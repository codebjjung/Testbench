module AXI_SLAVE;
	#(ADDR);
