module APB(
);
