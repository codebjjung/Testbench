module AXI_SLAVE;
	#(ADDR);
	endmodule
